`default_nettype none

//  Top level io for this module should stay the same to fit into the scan_wrapper.
//  The pin connections within the user_module are up to you,
//  although (if one is present) it is recommended to place a clock on io_in[0].
//  This allows use of the internal clock divider if you wish.
module user_module_341542971476279892(
  input [7:0] io_in, 
  output [7:0] io_out
);

  logo_341542971476279892 logo(
    .clk(io_in[0]),    
    .reset(io_in[1]),

    .img_sel(io_in[3:2]),
    .enable_horizontal(io_in[4]),

    .tx_out(io_out[0]),
    .h_sync(io_out[1]),
    .v_sync(io_out[2])
  );

endmodule

//  Any submodules should be included in this file,
//  so they are copied into the main TinyTapeout repo.
//  Appending your ID to any submodules you create 
//  ensures there are no clashes in full-chip simulation.

module logo_341542971476279892 (
    input clk,
    input reset,
    input [1:0] img_sel, //4 images
    input enable_horizontal, //enable lines
    
    output reg tx_out,
    output reg h_sync, //start of new line signal
    output reg v_sync  //start of new frame signal
  );

  reg       [9:0] rle_segment_counter;
  reg       [7:0] rle_pixel_counter;
  reg             rle_pixel_state;

  reg       [7:0] line_pixel_counter; //0 to IMG_WIDTH-1, pixels within a line

  reg       [9:0] next_rle_segment_counter;
  reg       [7:0] next_rle_pixel_counter;
  reg             next_rle_pixel_state;

  reg       [7:0] next_line_pixel_counter;

  reg       [7:0] current_rle_length; //length of current segment
  reg       [9:0] current_rle_n_segments; //number of segments in image
  
  reg             start_pixel;
  reg       [7:0] img_width; //max 255 with 8 bits

  //picture data
  parameter LEN_logoRLE = 111;
  parameter WIDTH_lambdaRLE = 41;
  parameter START_logoRLE = 1;
  wire [7:0] logoRLE [0:LEN_logoRLE-1];   //Edinburgh Hacklab logo
  
  parameter LEN_lambdaRLE = 207;
  parameter WIDTH_logoRLE = 41;
  parameter START_lambdaRLE = 1;
  wire [7:0] lambdaRLE [0:LEN_lambdaRLE-1]; //Lambda symbol

  parameter LEN_intRLE = 995;
  parameter WIDTH_intRLE = 125;
  parameter START_intRLE = 0;
  wire [7:0] intRLE [0:LEN_intRLE-1]; //lambda calculus diagram

  parameter LEN_amogusRLE = 301;
  parameter WIDTH_amogusRLE = 35;
  parameter START_amogusRLE = 1;
  wire [7:0] amogusRLE [0:LEN_amogusRLE-1]; //amogus meme

  assign logoRLE[0] = 41; assign logoRLE[1] = 136; assign logoRLE[2] = 5; assign logoRLE[3] = 35; assign logoRLE[4] = 7; assign logoRLE[5] = 33; assign logoRLE[6] = 8; assign logoRLE[7] = 33; assign logoRLE[8] = 9; assign logoRLE[9] = 32; assign logoRLE[10] = 2; assign logoRLE[11] = 3; assign logoRLE[12] = 4; assign logoRLE[13] = 32; assign logoRLE[14] = 2; assign logoRLE[15] = 4; assign logoRLE[16] = 3; assign logoRLE[17] = 31; assign logoRLE[18] = 2; assign logoRLE[19] = 6; assign logoRLE[20] = 3; assign logoRLE[21] = 30; assign logoRLE[22] = 2; assign logoRLE[23] = 6; assign logoRLE[24] = 3; assign logoRLE[25] = 38; assign logoRLE[26] = 3; assign logoRLE[27] = 39; assign logoRLE[28] = 2; assign logoRLE[29] = 39; assign logoRLE[30] = 3; assign logoRLE[31] = 37; assign logoRLE[32] = 4; assign logoRLE[33] = 37; assign logoRLE[34] = 4; assign logoRLE[35] = 36; assign logoRLE[36] = 5; assign logoRLE[37] = 36; assign logoRLE[38] = 6; assign logoRLE[39] = 35; assign logoRLE[40] = 6; assign logoRLE[41] = 34; assign logoRLE[42] = 7; assign logoRLE[43] = 34; assign logoRLE[44] = 7; assign logoRLE[45] = 33; assign logoRLE[46] = 5; assign logoRLE[47] = 1; assign logoRLE[48] = 2; assign logoRLE[49] = 33; assign logoRLE[50] = 5; assign logoRLE[51] = 1; assign logoRLE[52] = 3; assign logoRLE[53] = 31; assign logoRLE[54] = 6; assign logoRLE[55] = 1; assign logoRLE[56] = 3; assign logoRLE[57] = 31; assign logoRLE[58] = 5; assign logoRLE[59] = 2; assign logoRLE[60] = 3; assign logoRLE[61] = 30; assign logoRLE[62] = 6; assign logoRLE[63] = 2; assign logoRLE[64] = 3; assign logoRLE[65] = 30; assign logoRLE[66] = 5; assign logoRLE[67] = 4; assign logoRLE[68] = 3; assign logoRLE[69] = 28; assign logoRLE[70] = 6; assign logoRLE[71] = 4; assign logoRLE[72] = 3; assign logoRLE[73] = 5; assign logoRLE[74] = 2; assign logoRLE[75] = 21; assign logoRLE[76] = 5; assign logoRLE[77] = 5; assign logoRLE[78] = 3; assign logoRLE[79] = 5; assign logoRLE[80] = 2; assign logoRLE[81] = 20; assign logoRLE[82] = 6; assign logoRLE[83] = 5; assign logoRLE[84] = 4; assign logoRLE[85] = 4; assign logoRLE[86] = 2; assign logoRLE[87] = 20; assign logoRLE[88] = 5; assign logoRLE[89] = 7; assign logoRLE[90] = 4; assign logoRLE[91] = 2; assign logoRLE[92] = 3; assign logoRLE[93] = 20; assign logoRLE[94] = 5; assign logoRLE[95] = 7; assign logoRLE[96] = 9; assign logoRLE[97] = 19; assign logoRLE[98] = 6; assign logoRLE[99] = 7; assign logoRLE[100] = 8; assign logoRLE[101] = 20; assign logoRLE[102] = 5; assign logoRLE[103] = 9; assign logoRLE[104] = 7; assign logoRLE[105] = 20; assign logoRLE[106] = 5; assign logoRLE[107] = 10; assign logoRLE[108] = 5; assign logoRLE[109] = 175; assign logoRLE[110] = 41; 
  
  assign lambdaRLE[0] = 41; assign lambdaRLE[1] = 136; assign lambdaRLE[2] = 3; assign lambdaRLE[3] = 9; assign lambdaRLE[4] = 3; assign lambdaRLE[5] = 26; assign lambdaRLE[6] = 3; assign lambdaRLE[7] = 9; assign lambdaRLE[8] = 3; assign lambdaRLE[9] = 26; assign lambdaRLE[10] = 3; assign lambdaRLE[11] = 9; assign lambdaRLE[12] = 3; assign lambdaRLE[13] = 26; assign lambdaRLE[14] = 3; assign lambdaRLE[15] = 3; assign lambdaRLE[16] = 9; assign lambdaRLE[17] = 26; assign lambdaRLE[18] = 3; assign lambdaRLE[19] = 3; assign lambdaRLE[20] = 9; assign lambdaRLE[21] = 26; assign lambdaRLE[22] = 3; assign lambdaRLE[23] = 3; assign lambdaRLE[24] = 9; assign lambdaRLE[25] = 19; assign lambdaRLE[26] = 10; assign lambdaRLE[27] = 9; assign lambdaRLE[28] = 10; assign lambdaRLE[29] = 11; assign lambdaRLE[30] = 11; assign lambdaRLE[31] = 9; assign lambdaRLE[32] = 11; assign lambdaRLE[33] = 9; assign lambdaRLE[34] = 12; assign lambdaRLE[35] = 9; assign lambdaRLE[36] = 12; assign lambdaRLE[37] = 8; assign lambdaRLE[38] = 4; assign lambdaRLE[39] = 5; assign lambdaRLE[40] = 3; assign lambdaRLE[41] = 3; assign lambdaRLE[42] = 9; assign lambdaRLE[43] = 5; assign lambdaRLE[44] = 4; assign lambdaRLE[45] = 8; assign lambdaRLE[46] = 3; assign lambdaRLE[47] = 6; assign lambdaRLE[48] = 3; assign lambdaRLE[49] = 3; assign lambdaRLE[50] = 9; assign lambdaRLE[51] = 6; assign lambdaRLE[52] = 3; assign lambdaRLE[53] = 8; assign lambdaRLE[54] = 3; assign lambdaRLE[55] = 6; assign lambdaRLE[56] = 3; assign lambdaRLE[57] = 3; assign lambdaRLE[58] = 9; assign lambdaRLE[59] = 6; assign lambdaRLE[60] = 3; assign lambdaRLE[61] = 8; assign lambdaRLE[62] = 3; assign lambdaRLE[63] = 6; assign lambdaRLE[64] = 3; assign lambdaRLE[65] = 9; assign lambdaRLE[66] = 3; assign lambdaRLE[67] = 6; assign lambdaRLE[68] = 3; assign lambdaRLE[69] = 8; assign lambdaRLE[70] = 3; assign lambdaRLE[71] = 6; assign lambdaRLE[72] = 3; assign lambdaRLE[73] = 9; assign lambdaRLE[74] = 3; assign lambdaRLE[75] = 6; assign lambdaRLE[76] = 3; assign lambdaRLE[77] = 8; assign lambdaRLE[78] = 3; assign lambdaRLE[79] = 6; assign lambdaRLE[80] = 3; assign lambdaRLE[81] = 9; assign lambdaRLE[82] = 3; assign lambdaRLE[83] = 6; assign lambdaRLE[84] = 3; assign lambdaRLE[85] = 8; assign lambdaRLE[86] = 3; assign lambdaRLE[87] = 27; assign lambdaRLE[88] = 3; assign lambdaRLE[89] = 8; assign lambdaRLE[90] = 3; assign lambdaRLE[91] = 27; assign lambdaRLE[92] = 3; assign lambdaRLE[93] = 8; assign lambdaRLE[94] = 3; assign lambdaRLE[95] = 27; assign lambdaRLE[96] = 3; assign lambdaRLE[97] = 8; assign lambdaRLE[98] = 3; assign lambdaRLE[99] = 6; assign lambdaRLE[100] = 3; assign lambdaRLE[101] = 3; assign lambdaRLE[102] = 3; assign lambdaRLE[103] = 3; assign lambdaRLE[104] = 3; assign lambdaRLE[105] = 6; assign lambdaRLE[106] = 3; assign lambdaRLE[107] = 8; assign lambdaRLE[108] = 3; assign lambdaRLE[109] = 6; assign lambdaRLE[110] = 3; assign lambdaRLE[111] = 3; assign lambdaRLE[112] = 3; assign lambdaRLE[113] = 3; assign lambdaRLE[114] = 3; assign lambdaRLE[115] = 6; assign lambdaRLE[116] = 3; assign lambdaRLE[117] = 8; assign lambdaRLE[118] = 3; assign lambdaRLE[119] = 6; assign lambdaRLE[120] = 3; assign lambdaRLE[121] = 3; assign lambdaRLE[122] = 3; assign lambdaRLE[123] = 3; assign lambdaRLE[124] = 3; assign lambdaRLE[125] = 6; assign lambdaRLE[126] = 3; assign lambdaRLE[127] = 8; assign lambdaRLE[128] = 3; assign lambdaRLE[129] = 6; assign lambdaRLE[130] = 3; assign lambdaRLE[131] = 3; assign lambdaRLE[132] = 3; assign lambdaRLE[133] = 3; assign lambdaRLE[134] = 3; assign lambdaRLE[135] = 6; assign lambdaRLE[136] = 3; assign lambdaRLE[137] = 8; assign lambdaRLE[138] = 3; assign lambdaRLE[139] = 6; assign lambdaRLE[140] = 3; assign lambdaRLE[141] = 3; assign lambdaRLE[142] = 3; assign lambdaRLE[143] = 3; assign lambdaRLE[144] = 3; assign lambdaRLE[145] = 6; assign lambdaRLE[146] = 3; assign lambdaRLE[147] = 8; assign lambdaRLE[148] = 4; assign lambdaRLE[149] = 5; assign lambdaRLE[150] = 3; assign lambdaRLE[151] = 3; assign lambdaRLE[152] = 3; assign lambdaRLE[153] = 3; assign lambdaRLE[154] = 3; assign lambdaRLE[155] = 5; assign lambdaRLE[156] = 4; assign lambdaRLE[157] = 8; assign lambdaRLE[158] = 12; assign lambdaRLE[159] = 9; assign lambdaRLE[160] = 12; assign lambdaRLE[161] = 9; assign lambdaRLE[162] = 11; assign lambdaRLE[163] = 9; assign lambdaRLE[164] = 11; assign lambdaRLE[165] = 11; assign lambdaRLE[166] = 10; assign lambdaRLE[167] = 9; assign lambdaRLE[168] = 10; assign lambdaRLE[169] = 19; assign lambdaRLE[170] = 3; assign lambdaRLE[171] = 3; assign lambdaRLE[172] = 3; assign lambdaRLE[173] = 3; assign lambdaRLE[174] = 3; assign lambdaRLE[175] = 26; assign lambdaRLE[176] = 3; assign lambdaRLE[177] = 3; assign lambdaRLE[178] = 3; assign lambdaRLE[179] = 3; assign lambdaRLE[180] = 3; assign lambdaRLE[181] = 26; assign lambdaRLE[182] = 3; assign lambdaRLE[183] = 3; assign lambdaRLE[184] = 3; assign lambdaRLE[185] = 3; assign lambdaRLE[186] = 3; assign lambdaRLE[187] = 26; assign lambdaRLE[188] = 3; assign lambdaRLE[189] = 3; assign lambdaRLE[190] = 3; assign lambdaRLE[191] = 3; assign lambdaRLE[192] = 3; assign lambdaRLE[193] = 26; assign lambdaRLE[194] = 3; assign lambdaRLE[195] = 3; assign lambdaRLE[196] = 3; assign lambdaRLE[197] = 3; assign lambdaRLE[198] = 3; assign lambdaRLE[199] = 26; assign lambdaRLE[200] = 3; assign lambdaRLE[201] = 3; assign lambdaRLE[202] = 3; assign lambdaRLE[203] = 3; assign lambdaRLE[204] = 3; assign lambdaRLE[205] = 136; assign lambdaRLE[206] = 41;

  assign intRLE[0] = 126; assign intRLE[1] = 7; assign intRLE[2] = 1; assign intRLE[3] = 115; assign intRLE[4] = 3; assign intRLE[5] = 1; assign intRLE[6] = 3; assign intRLE[7] = 1; assign intRLE[8] = 107; assign intRLE[9] = 1; assign intRLE[10] = 3; assign intRLE[11] = 1; assign intRLE[12] = 8; assign intRLE[13] = 5; assign intRLE[14] = 2; assign intRLE[15] = 115; assign intRLE[16] = 7; assign intRLE[17] = 1; assign intRLE[18] = 107; assign intRLE[19] = 1; assign intRLE[20] = 3; assign intRLE[21] = 1; assign intRLE[22] = 3; assign intRLE[23] = 1; assign intRLE[24] = 8; assign intRLE[25] = 1; assign intRLE[26] = 2; assign intRLE[27] = 115; assign intRLE[28] = 7; assign intRLE[29] = 1; assign intRLE[30] = 3; assign intRLE[31] = 1; assign intRLE[32] = 103; assign intRLE[33] = 1; assign intRLE[34] = 3; assign intRLE[35] = 1; assign intRLE[36] = 3; assign intRLE[37] = 1; assign intRLE[38] = 8; assign intRLE[39] = 1; assign intRLE[40] = 3; assign intRLE[41] = 1; assign intRLE[42] = 2; assign intRLE[43] = 99; assign intRLE[44] = 2; assign intRLE[45] = 5; assign intRLE[46] = 3; assign intRLE[47] = 1; assign intRLE[48] = 8; assign intRLE[49] = 1; assign intRLE[50] = 3; assign intRLE[51] = 1; assign intRLE[52] = 7; assign intRLE[53] = 1; assign intRLE[54] = 95; assign intRLE[55] = 1; assign intRLE[56] = 7; assign intRLE[57] = 1; assign intRLE[58] = 8; assign intRLE[59] = 1; assign intRLE[60] = 3; assign intRLE[61] = 1; assign intRLE[62] = 2; assign intRLE[63] = 99; assign intRLE[64] = 2; assign intRLE[65] = 1; assign intRLE[66] = 7; assign intRLE[67] = 1; assign intRLE[68] = 8; assign intRLE[69] = 1; assign intRLE[70] = 3; assign intRLE[71] = 1; assign intRLE[72] = 3; assign intRLE[73] = 1; assign intRLE[74] = 3; assign intRLE[75] = 1; assign intRLE[76] = 91; assign intRLE[77] = 1; assign intRLE[78] = 3; assign intRLE[79] = 1; assign intRLE[80] = 7; assign intRLE[81] = 1; assign intRLE[82] = 8; assign intRLE[83] = 1; assign intRLE[84] = 3; assign intRLE[85] = 1; assign intRLE[86] = 2; assign intRLE[87] = 99; assign intRLE[88] = 2; assign intRLE[89] = 1; assign intRLE[90] = 7; assign intRLE[91] = 1; assign intRLE[92] = 8; assign intRLE[93] = 1; assign intRLE[94] = 3; assign intRLE[95] = 1; assign intRLE[96] = 3; assign intRLE[97] = 1; assign intRLE[98] = 3; assign intRLE[99] = 1; assign intRLE[100] = 3; assign intRLE[101] = 1; assign intRLE[102] = 27; assign intRLE[103] = 1; assign intRLE[104] = 39; assign intRLE[105] = 1; assign intRLE[106] = 19; assign intRLE[107] = 1; assign intRLE[108] = 3; assign intRLE[109] = 1; assign intRLE[110] = 7; assign intRLE[111] = 1; assign intRLE[112] = 8; assign intRLE[113] = 1; assign intRLE[114] = 3; assign intRLE[115] = 1; assign intRLE[116] = 2; assign intRLE[117] = 99; assign intRLE[118] = 2; assign intRLE[119] = 1; assign intRLE[120] = 7; assign intRLE[121] = 1; assign intRLE[122] = 8; assign intRLE[123] = 1; assign intRLE[124] = 3; assign intRLE[125] = 1; assign intRLE[126] = 3; assign intRLE[127] = 1; assign intRLE[128] = 3; assign intRLE[129] = 1; assign intRLE[130] = 3; assign intRLE[131] = 1; assign intRLE[132] = 7; assign intRLE[133] = 1; assign intRLE[134] = 19; assign intRLE[135] = 1; assign intRLE[136] = 3; assign intRLE[137] = 1; assign intRLE[138] = 23; assign intRLE[139] = 1; assign intRLE[140] = 11; assign intRLE[141] = 1; assign intRLE[142] = 3; assign intRLE[143] = 1; assign intRLE[144] = 15; assign intRLE[145] = 1; assign intRLE[146] = 3; assign intRLE[147] = 1; assign intRLE[148] = 7; assign intRLE[149] = 1; assign intRLE[150] = 8; assign intRLE[151] = 1; assign intRLE[152] = 3; assign intRLE[153] = 1; assign intRLE[154] = 3; assign intRLE[155] = 1; assign intRLE[156] = 2; assign intRLE[157] = 95; assign intRLE[158] = 2; assign intRLE[159] = 1; assign intRLE[160] = 7; assign intRLE[161] = 1; assign intRLE[162] = 8; assign intRLE[163] = 1; assign intRLE[164] = 3; assign intRLE[165] = 1; assign intRLE[166] = 3; assign intRLE[167] = 1; assign intRLE[168] = 3; assign intRLE[169] = 1; assign intRLE[170] = 3; assign intRLE[171] = 1; assign intRLE[172] = 3; assign intRLE[173] = 1; assign intRLE[174] = 3; assign intRLE[175] = 1; assign intRLE[176] = 19; assign intRLE[177] = 1; assign intRLE[178] = 3; assign intRLE[179] = 1; assign intRLE[180] = 19; assign intRLE[181] = 1; assign intRLE[182] = 3; assign intRLE[183] = 1; assign intRLE[184] = 7; assign intRLE[185] = 1; assign intRLE[186] = 3; assign intRLE[187] = 1; assign intRLE[188] = 3; assign intRLE[189] = 1; assign intRLE[190] = 11; assign intRLE[191] = 1; assign intRLE[192] = 3; assign intRLE[193] = 1; assign intRLE[194] = 3; assign intRLE[195] = 1; assign intRLE[196] = 7; assign intRLE[197] = 1; assign intRLE[198] = 8; assign intRLE[199] = 1; assign intRLE[200] = 3; assign intRLE[201] = 1; assign intRLE[202] = 3; assign intRLE[203] = 1; assign intRLE[204] = 3; assign intRLE[205] = 1; assign intRLE[206] = 3; assign intRLE[207] = 1; assign intRLE[208] = 2; assign intRLE[209] = 47; assign intRLE[210] = 2; assign intRLE[211] = 1; assign intRLE[212] = 3; assign intRLE[213] = 1; assign intRLE[214] = 2; assign intRLE[215] = 7; assign intRLE[216] = 1; assign intRLE[217] = 23; assign intRLE[218] = 2; assign intRLE[219] = 1; assign intRLE[220] = 7; assign intRLE[221] = 1; assign intRLE[222] = 8; assign intRLE[223] = 1; assign intRLE[224] = 3; assign intRLE[225] = 1; assign intRLE[226] = 3; assign intRLE[227] = 1; assign intRLE[228] = 3; assign intRLE[229] = 1; assign intRLE[230] = 3; assign intRLE[231] = 1; assign intRLE[232] = 3; assign intRLE[233] = 1; assign intRLE[234] = 3; assign intRLE[235] = 1; assign intRLE[236] = 3; assign intRLE[237] = 1; assign intRLE[238] = 15; assign intRLE[239] = 1; assign intRLE[240] = 3; assign intRLE[241] = 1; assign intRLE[242] = 3; assign intRLE[243] = 1; assign intRLE[244] = 15; assign intRLE[245] = 1; assign intRLE[246] = 3; assign intRLE[247] = 1; assign intRLE[248] = 3; assign intRLE[249] = 1; assign intRLE[250] = 3; assign intRLE[251] = 1; assign intRLE[252] = 3; assign intRLE[253] = 1; assign intRLE[254] = 3; assign intRLE[255] = 1; assign intRLE[256] = 11; assign intRLE[257] = 1; assign intRLE[258] = 3; assign intRLE[259] = 1; assign intRLE[260] = 3; assign intRLE[261] = 1; assign intRLE[262] = 7; assign intRLE[263] = 1; assign intRLE[264] = 8; assign intRLE[265] = 1; assign intRLE[266] = 3; assign intRLE[267] = 1; assign intRLE[268] = 3; assign intRLE[269] = 1; assign intRLE[270] = 3; assign intRLE[271] = 1; assign intRLE[272] = 3; assign intRLE[273] = 1; assign intRLE[274] = 3; assign intRLE[275] = 1; assign intRLE[276] = 3; assign intRLE[277] = 1; assign intRLE[278] = 2; assign intRLE[279] = 15; assign intRLE[280] = 2; assign intRLE[281] = 1; assign intRLE[282] = 2; assign intRLE[283] = 19; assign intRLE[284] = 2; assign intRLE[285] = 1; assign intRLE[286] = 3; assign intRLE[287] = 1; assign intRLE[288] = 3; assign intRLE[289] = 5; assign intRLE[290] = 3; assign intRLE[291] = 1; assign intRLE[292] = 2; assign intRLE[293] = 15; assign intRLE[294] = 2; assign intRLE[295] = 1; assign intRLE[296] = 3; assign intRLE[297] = 1; assign intRLE[298] = 7; assign intRLE[299] = 1; assign intRLE[300] = 8; assign intRLE[301] = 1; assign intRLE[302] = 3; assign intRLE[303] = 1; assign intRLE[304] = 3; assign intRLE[305] = 1; assign intRLE[306] = 3; assign intRLE[307] = 1; assign intRLE[308] = 3; assign intRLE[309] = 1; assign intRLE[310] = 3; assign intRLE[311] = 1; assign intRLE[312] = 3; assign intRLE[313] = 1; assign intRLE[314] = 3; assign intRLE[315] = 1; assign intRLE[316] = 11; assign intRLE[317] = 1; assign intRLE[318] = 3; assign intRLE[319] = 1; assign intRLE[320] = 3; assign intRLE[321] = 1; assign intRLE[322] = 3; assign intRLE[323] = 1; assign intRLE[324] = 7; assign intRLE[325] = 1; assign intRLE[326] = 7; assign intRLE[327] = 1; assign intRLE[328] = 3; assign intRLE[329] = 1; assign intRLE[330] = 3; assign intRLE[331] = 1; assign intRLE[332] = 7; assign intRLE[333] = 1; assign intRLE[334] = 3; assign intRLE[335] = 1; assign intRLE[336] = 3; assign intRLE[337] = 1; assign intRLE[338] = 7; assign intRLE[339] = 1; assign intRLE[340] = 3; assign intRLE[341] = 1; assign intRLE[342] = 3; assign intRLE[343] = 1; assign intRLE[344] = 7; assign intRLE[345] = 1; assign intRLE[346] = 8; assign intRLE[347] = 1; assign intRLE[348] = 3; assign intRLE[349] = 1; assign intRLE[350] = 3; assign intRLE[351] = 1; assign intRLE[352] = 3; assign intRLE[353] = 1; assign intRLE[354] = 3; assign intRLE[355] = 1; assign intRLE[356] = 3; assign intRLE[357] = 1; assign intRLE[358] = 3; assign intRLE[359] = 1; assign intRLE[360] = 2; assign intRLE[361] = 15; assign intRLE[362] = 2; assign intRLE[363] = 1; assign intRLE[364] = 3; assign intRLE[365] = 1; assign intRLE[366] = 2; assign intRLE[367] = 15; assign intRLE[368] = 2; assign intRLE[369] = 1; assign intRLE[370] = 3; assign intRLE[371] = 5; assign intRLE[372] = 7; assign intRLE[373] = 1; assign intRLE[374] = 3; assign intRLE[375] = 1; assign intRLE[376] = 2; assign intRLE[377] = 11; assign intRLE[378] = 2; assign intRLE[379] = 1; assign intRLE[380] = 3; assign intRLE[381] = 1; assign intRLE[382] = 7; assign intRLE[383] = 1; assign intRLE[384] = 8; assign intRLE[385] = 1; assign intRLE[386] = 3; assign intRLE[387] = 1; assign intRLE[388] = 3; assign intRLE[389] = 1; assign intRLE[390] = 3; assign intRLE[391] = 1; assign intRLE[392] = 3; assign intRLE[393] = 1; assign intRLE[394] = 3; assign intRLE[395] = 1; assign intRLE[396] = 3; assign intRLE[397] = 1; assign intRLE[398] = 3; assign intRLE[399] = 1; assign intRLE[400] = 7; assign intRLE[401] = 1; assign intRLE[402] = 3; assign intRLE[403] = 1; assign intRLE[404] = 3; assign intRLE[405] = 1; assign intRLE[406] = 3; assign intRLE[407] = 1; assign intRLE[408] = 3; assign intRLE[409] = 1; assign intRLE[410] = 3; assign intRLE[411] = 1; assign intRLE[412] = 3; assign intRLE[413] = 1; assign intRLE[414] = 3; assign intRLE[415] = 1; assign intRLE[416] = 3; assign intRLE[417] = 1; assign intRLE[418] = 3; assign intRLE[419] = 1; assign intRLE[420] = 11; assign intRLE[421] = 1; assign intRLE[422] = 3; assign intRLE[423] = 1; assign intRLE[424] = 3; assign intRLE[425] = 1; assign intRLE[426] = 3; assign intRLE[427] = 1; assign intRLE[428] = 3; assign intRLE[429] = 1; assign intRLE[430] = 3; assign intRLE[431] = 1; assign intRLE[432] = 3; assign intRLE[433] = 1; assign intRLE[434] = 7; assign intRLE[435] = 1; assign intRLE[436] = 8; assign intRLE[437] = 1; assign intRLE[438] = 3; assign intRLE[439] = 1; assign intRLE[440] = 3; assign intRLE[441] = 1; assign intRLE[442] = 3; assign intRLE[443] = 1; assign intRLE[444] = 3; assign intRLE[445] = 1; assign intRLE[446] = 3; assign intRLE[447] = 1; assign intRLE[448] = 3; assign intRLE[449] = 1; assign intRLE[450] = 3; assign intRLE[451] = 1; assign intRLE[452] = 2; assign intRLE[453] = 11; assign intRLE[454] = 2; assign intRLE[455] = 1; assign intRLE[456] = 3; assign intRLE[457] = 1; assign intRLE[458] = 3; assign intRLE[459] = 5; assign intRLE[460] = 3; assign intRLE[461] = 5; assign intRLE[462] = 3; assign intRLE[463] = 5; assign intRLE[464] = 11; assign intRLE[465] = 1; assign intRLE[466] = 3; assign intRLE[467] = 1; assign intRLE[468] = 3; assign intRLE[469] = 1; assign intRLE[470] = 3; assign intRLE[471] = 5; assign intRLE[472] = 3; assign intRLE[473] = 1; assign intRLE[474] = 3; assign intRLE[475] = 1; assign intRLE[476] = 7; assign intRLE[477] = 1; assign intRLE[478] = 8; assign intRLE[479] = 1; assign intRLE[480] = 3; assign intRLE[481] = 1; assign intRLE[482] = 3; assign intRLE[483] = 1; assign intRLE[484] = 3; assign intRLE[485] = 1; assign intRLE[486] = 3; assign intRLE[487] = 1; assign intRLE[488] = 3; assign intRLE[489] = 1; assign intRLE[490] = 3; assign intRLE[491] = 1; assign intRLE[492] = 3; assign intRLE[493] = 1; assign intRLE[494] = 3; assign intRLE[495] = 1; assign intRLE[496] = 3; assign intRLE[497] = 1; assign intRLE[498] = 3; assign intRLE[499] = 1; assign intRLE[500] = 3; assign intRLE[501] = 1; assign intRLE[502] = 3; assign intRLE[503] = 1; assign intRLE[504] = 7; assign intRLE[505] = 1; assign intRLE[506] = 3; assign intRLE[507] = 1; assign intRLE[508] = 11; assign intRLE[509] = 1; assign intRLE[510] = 11; assign intRLE[511] = 1; assign intRLE[512] = 3; assign intRLE[513] = 1; assign intRLE[514] = 3; assign intRLE[515] = 1; assign intRLE[516] = 3; assign intRLE[517] = 1; assign intRLE[518] = 7; assign intRLE[519] = 1; assign intRLE[520] = 3; assign intRLE[521] = 1; assign intRLE[522] = 7; assign intRLE[523] = 1; assign intRLE[524] = 8; assign intRLE[525] = 1; assign intRLE[526] = 3; assign intRLE[527] = 1; assign intRLE[528] = 3; assign intRLE[529] = 1; assign intRLE[530] = 3; assign intRLE[531] = 1; assign intRLE[532] = 3; assign intRLE[533] = 1; assign intRLE[534] = 3; assign intRLE[535] = 1; assign intRLE[536] = 3; assign intRLE[537] = 1; assign intRLE[538] = 3; assign intRLE[539] = 1; assign intRLE[540] = 3; assign intRLE[541] = 5; assign intRLE[542] = 3; assign intRLE[543] = 1; assign intRLE[544] = 3; assign intRLE[545] = 1; assign intRLE[546] = 3; assign intRLE[547] = 1; assign intRLE[548] = 7; assign intRLE[549] = 5; assign intRLE[550] = 11; assign intRLE[551] = 1; assign intRLE[552] = 11; assign intRLE[553] = 1; assign intRLE[554] = 3; assign intRLE[555] = 1; assign intRLE[556] = 3; assign intRLE[557] = 5; assign intRLE[558] = 7; assign intRLE[559] = 1; assign intRLE[560] = 3; assign intRLE[561] = 1; assign intRLE[562] = 7; assign intRLE[563] = 1; assign intRLE[564] = 8; assign intRLE[565] = 1; assign intRLE[566] = 3; assign intRLE[567] = 1; assign intRLE[568] = 3; assign intRLE[569] = 1; assign intRLE[570] = 3; assign intRLE[571] = 1; assign intRLE[572] = 3; assign intRLE[573] = 1; assign intRLE[574] = 3; assign intRLE[575] = 1; assign intRLE[576] = 3; assign intRLE[577] = 1; assign intRLE[578] = 3; assign intRLE[579] = 1; assign intRLE[580] = 7; assign intRLE[581] = 1; assign intRLE[582] = 3; assign intRLE[583] = 1; assign intRLE[584] = 3; assign intRLE[585] = 1; assign intRLE[586] = 3; assign intRLE[587] = 1; assign intRLE[588] = 7; assign intRLE[589] = 1; assign intRLE[590] = 15; assign intRLE[591] = 1; assign intRLE[592] = 11; assign intRLE[593] = 1; assign intRLE[594] = 3; assign intRLE[595] = 1; assign intRLE[596] = 3; assign intRLE[597] = 1; assign intRLE[598] = 11; assign intRLE[599] = 1; assign intRLE[600] = 3; assign intRLE[601] = 1; assign intRLE[602] = 7; assign intRLE[603] = 1; assign intRLE[604] = 8; assign intRLE[605] = 1; assign intRLE[606] = 3; assign intRLE[607] = 1; assign intRLE[608] = 3; assign intRLE[609] = 1; assign intRLE[610] = 3; assign intRLE[611] = 1; assign intRLE[612] = 3; assign intRLE[613] = 1; assign intRLE[614] = 3; assign intRLE[615] = 1; assign intRLE[616] = 3; assign intRLE[617] = 1; assign intRLE[618] = 3; assign intRLE[619] = 1; assign intRLE[620] = 7; assign intRLE[621] = 5; assign intRLE[622] = 3; assign intRLE[623] = 1; assign intRLE[624] = 3; assign intRLE[625] = 9; assign intRLE[626] = 15; assign intRLE[627] = 1; assign intRLE[628] = 11; assign intRLE[629] = 1; assign intRLE[630] = 3; assign intRLE[631] = 5; assign intRLE[632] = 11; assign intRLE[633] = 1; assign intRLE[634] = 3; assign intRLE[635] = 1; assign intRLE[636] = 7; assign intRLE[637] = 1; assign intRLE[638] = 8; assign intRLE[639] = 1; assign intRLE[640] = 3; assign intRLE[641] = 1; assign intRLE[642] = 3; assign intRLE[643] = 1; assign intRLE[644] = 3; assign intRLE[645] = 1; assign intRLE[646] = 3; assign intRLE[647] = 1; assign intRLE[648] = 3; assign intRLE[649] = 1; assign intRLE[650] = 3; assign intRLE[651] = 1; assign intRLE[652] = 3; assign intRLE[653] = 1; assign intRLE[654] = 7; assign intRLE[655] = 1; assign intRLE[656] = 7; assign intRLE[657] = 1; assign intRLE[658] = 3; assign intRLE[659] = 1; assign intRLE[660] = 23; assign intRLE[661] = 1; assign intRLE[662] = 11; assign intRLE[663] = 1; assign intRLE[664] = 3; assign intRLE[665] = 1; assign intRLE[666] = 15; assign intRLE[667] = 1; assign intRLE[668] = 3; assign intRLE[669] = 1; assign intRLE[670] = 7; assign intRLE[671] = 1; assign intRLE[672] = 8; assign intRLE[673] = 1; assign intRLE[674] = 3; assign intRLE[675] = 1; assign intRLE[676] = 3; assign intRLE[677] = 1; assign intRLE[678] = 3; assign intRLE[679] = 1; assign intRLE[680] = 3; assign intRLE[681] = 1; assign intRLE[682] = 3; assign intRLE[683] = 1; assign intRLE[684] = 3; assign intRLE[685] = 1; assign intRLE[686] = 3; assign intRLE[687] = 9; assign intRLE[688] = 7; assign intRLE[689] = 5; assign intRLE[690] = 23; assign intRLE[691] = 1; assign intRLE[692] = 11; assign intRLE[693] = 5; assign intRLE[694] = 15; assign intRLE[695] = 1; assign intRLE[696] = 3; assign intRLE[697] = 1; assign intRLE[698] = 7; assign intRLE[699] = 1; assign intRLE[700] = 8; assign intRLE[701] = 1; assign intRLE[702] = 3; assign intRLE[703] = 1; assign intRLE[704] = 3; assign intRLE[705] = 1; assign intRLE[706] = 3; assign intRLE[707] = 1; assign intRLE[708] = 3; assign intRLE[709] = 1; assign intRLE[710] = 3; assign intRLE[711] = 1; assign intRLE[712] = 3; assign intRLE[713] = 1; assign intRLE[714] = 3; assign intRLE[715] = 1; assign intRLE[716] = 15; assign intRLE[717] = 1; assign intRLE[718] = 27; assign intRLE[719] = 1; assign intRLE[720] = 15; assign intRLE[721] = 1; assign intRLE[722] = 15; assign intRLE[723] = 1; assign intRLE[724] = 3; assign intRLE[725] = 1; assign intRLE[726] = 7; assign intRLE[727] = 1; assign intRLE[728] = 8; assign intRLE[729] = 1; assign intRLE[730] = 3; assign intRLE[731] = 1; assign intRLE[732] = 3; assign intRLE[733] = 1; assign intRLE[734] = 3; assign intRLE[735] = 1; assign intRLE[736] = 3; assign intRLE[737] = 1; assign intRLE[738] = 3; assign intRLE[739] = 1; assign intRLE[740] = 3; assign intRLE[741] = 5; assign intRLE[742] = 15; assign intRLE[743] = 1; assign intRLE[744] = 27; assign intRLE[745] = 1; assign intRLE[746] = 15; assign intRLE[747] = 17; assign intRLE[748] = 3; assign intRLE[749] = 1; assign intRLE[750] = 7; assign intRLE[751] = 1; assign intRLE[752] = 8; assign intRLE[753] = 1; assign intRLE[754] = 3; assign intRLE[755] = 1; assign intRLE[756] = 3; assign intRLE[757] = 1; assign intRLE[758] = 3; assign intRLE[759] = 1; assign intRLE[760] = 3; assign intRLE[761] = 1; assign intRLE[762] = 3; assign intRLE[763] = 1; assign intRLE[764] = 3; assign intRLE[765] = 1; assign intRLE[766] = 19; assign intRLE[767] = 1; assign intRLE[768] = 27; assign intRLE[769] = 1; assign intRLE[770] = 15; assign intRLE[771] = 1; assign intRLE[772] = 19; assign intRLE[773] = 1; assign intRLE[774] = 7; assign intRLE[775] = 1; assign intRLE[776] = 8; assign intRLE[777] = 1; assign intRLE[778] = 3; assign intRLE[779] = 1; assign intRLE[780] = 3; assign intRLE[781] = 1; assign intRLE[782] = 3; assign intRLE[783] = 1; assign intRLE[784] = 3; assign intRLE[785] = 1; assign intRLE[786] = 3; assign intRLE[787] = 5; assign intRLE[788] = 19; assign intRLE[789] = 1; assign intRLE[790] = 27; assign intRLE[791] = 17; assign intRLE[792] = 19; assign intRLE[793] = 1; assign intRLE[794] = 7; assign intRLE[795] = 1; assign intRLE[796] = 8; assign intRLE[797] = 1; assign intRLE[798] = 3; assign intRLE[799] = 1; assign intRLE[800] = 3; assign intRLE[801] = 1; assign intRLE[802] = 3; assign intRLE[803] = 1; assign intRLE[804] = 3; assign intRLE[805] = 1; assign intRLE[806] = 7; assign intRLE[807] = 1; assign intRLE[808] = 19; assign intRLE[809] = 1; assign intRLE[810] = 27; assign intRLE[811] = 1; assign intRLE[812] = 35; assign intRLE[813] = 1; assign intRLE[814] = 7; assign intRLE[815] = 1; assign intRLE[816] = 8; assign intRLE[817] = 1; assign intRLE[818] = 3; assign intRLE[819] = 1; assign intRLE[820] = 3; assign intRLE[821] = 1; assign intRLE[822] = 3; assign intRLE[823] = 1; assign intRLE[824] = 3; assign intRLE[825] = 1; assign intRLE[826] = 7; assign intRLE[827] = 21; assign intRLE[828] = 27; assign intRLE[829] = 1; assign intRLE[830] = 35; assign intRLE[831] = 1; assign intRLE[832] = 7; assign intRLE[833] = 1; assign intRLE[834] = 8; assign intRLE[835] = 1; assign intRLE[836] = 3; assign intRLE[837] = 1; assign intRLE[838] = 3; assign intRLE[839] = 1; assign intRLE[840] = 3; assign intRLE[841] = 1; assign intRLE[842] = 3; assign intRLE[843] = 1; assign intRLE[844] = 7; assign intRLE[845] = 1; assign intRLE[846] = 47; assign intRLE[847] = 1; assign intRLE[848] = 35; assign intRLE[849] = 1; assign intRLE[850] = 7; assign intRLE[851] = 1; assign intRLE[852] = 8; assign intRLE[853] = 1; assign intRLE[854] = 3; assign intRLE[855] = 1; assign intRLE[856] = 3; assign intRLE[857] = 1; assign intRLE[858] = 3; assign intRLE[859] = 1; assign intRLE[860] = 3; assign intRLE[861] = 9; assign intRLE[862] = 47; assign intRLE[863] = 1; assign intRLE[864] = 35; assign intRLE[865] = 1; assign intRLE[866] = 7; assign intRLE[867] = 1; assign intRLE[868] = 8; assign intRLE[869] = 1; assign intRLE[870] = 3; assign intRLE[871] = 1; assign intRLE[872] = 3; assign intRLE[873] = 1; assign intRLE[874] = 3; assign intRLE[875] = 1; assign intRLE[876] = 3; assign intRLE[877] = 1; assign intRLE[878] = 55; assign intRLE[879] = 1; assign intRLE[880] = 35; assign intRLE[881] = 1; assign intRLE[882] = 7; assign intRLE[883] = 1; assign intRLE[884] = 8; assign intRLE[885] = 1; assign intRLE[886] = 3; assign intRLE[887] = 1; assign intRLE[888] = 3; assign intRLE[889] = 1; assign intRLE[890] = 3; assign intRLE[891] = 5; assign intRLE[892] = 55; assign intRLE[893] = 1; assign intRLE[894] = 35; assign intRLE[895] = 1; assign intRLE[896] = 7; assign intRLE[897] = 1; assign intRLE[898] = 8; assign intRLE[899] = 1; assign intRLE[900] = 3; assign intRLE[901] = 1; assign intRLE[902] = 3; assign intRLE[903] = 1; assign intRLE[904] = 7; assign intRLE[905] = 1; assign intRLE[906] = 55; assign intRLE[907] = 1; assign intRLE[908] = 35; assign intRLE[909] = 1; assign intRLE[910] = 7; assign intRLE[911] = 1; assign intRLE[912] = 8; assign intRLE[913] = 1; assign intRLE[914] = 3; assign intRLE[915] = 1; assign intRLE[916] = 3; assign intRLE[917] = 1; assign intRLE[918] = 7; assign intRLE[919] = 57; assign intRLE[920] = 35; assign intRLE[921] = 1; assign intRLE[922] = 7; assign intRLE[923] = 1; assign intRLE[924] = 8; assign intRLE[925] = 1; assign intRLE[926] = 3; assign intRLE[927] = 1; assign intRLE[928] = 3; assign intRLE[929] = 1; assign intRLE[930] = 7; assign intRLE[931] = 1; assign intRLE[932] = 91; assign intRLE[933] = 1; assign intRLE[934] = 7; assign intRLE[935] = 1; assign intRLE[936] = 8; assign intRLE[937] = 1; assign intRLE[938] = 3; assign intRLE[939] = 1; assign intRLE[940] = 3; assign intRLE[941] = 9; assign intRLE[942] = 91; assign intRLE[943] = 1; assign intRLE[944] = 7; assign intRLE[945] = 1; assign intRLE[946] = 8; assign intRLE[947] = 1; assign intRLE[948] = 3; assign intRLE[949] = 1; assign intRLE[950] = 3; assign intRLE[951] = 1; assign intRLE[952] = 99; assign intRLE[953] = 1; assign intRLE[954] = 7; assign intRLE[955] = 1; assign intRLE[956] = 8; assign intRLE[957] = 1; assign intRLE[958] = 3; assign intRLE[959] = 5; assign intRLE[960] = 99; assign intRLE[961] = 1; assign intRLE[962] = 7; assign intRLE[963] = 1; assign intRLE[964] = 8; assign intRLE[965] = 1; assign intRLE[966] = 7; assign intRLE[967] = 1; assign intRLE[968] = 99; assign intRLE[969] = 1; assign intRLE[970] = 7; assign intRLE[971] = 1; assign intRLE[972] = 8; assign intRLE[973] = 1; assign intRLE[974] = 7; assign intRLE[975] = 101; assign intRLE[976] = 7; assign intRLE[977] = 1; assign intRLE[978] = 8; assign intRLE[979] = 1; assign intRLE[980] = 107; assign intRLE[981] = 1; assign intRLE[982] = 7; assign intRLE[983] = 1; assign intRLE[984] = 8; assign intRLE[985] = 1; assign intRLE[986] = 107; assign intRLE[987] = 9; assign intRLE[988] = 8; assign intRLE[989] = 1; assign intRLE[990] = 107; assign intRLE[991] = 1; assign intRLE[992] = 16; assign intRLE[993] = 109; assign intRLE[994] = 135;

  assign amogusRLE[0] = 35; assign amogusRLE[1] = 75; assign amogusRLE[2] = 1; assign amogusRLE[3] = 3; assign amogusRLE[4] = 1; assign amogusRLE[5] = 1; assign amogusRLE[6] = 1; assign amogusRLE[7] = 3; assign amogusRLE[8] = 1; assign amogusRLE[9] = 3; assign amogusRLE[10] = 2; assign amogusRLE[11] = 2; assign amogusRLE[12] = 1; assign amogusRLE[13] = 1; assign amogusRLE[14] = 1; assign amogusRLE[15] = 1; assign amogusRLE[16] = 3; assign amogusRLE[17] = 9; assign amogusRLE[18] = 1; assign amogusRLE[19] = 1; assign amogusRLE[20] = 1; assign amogusRLE[21] = 1; assign amogusRLE[22] = 1; assign amogusRLE[23] = 1; assign amogusRLE[24] = 1; assign amogusRLE[25] = 1; assign amogusRLE[26] = 1; assign amogusRLE[27] = 1; assign amogusRLE[28] = 1; assign amogusRLE[29] = 1; assign amogusRLE[30] = 1; assign amogusRLE[31] = 1; assign amogusRLE[32] = 1; assign amogusRLE[33] = 4; assign amogusRLE[34] = 1; assign amogusRLE[35] = 1; assign amogusRLE[36] = 1; assign amogusRLE[37] = 1; assign amogusRLE[38] = 1; assign amogusRLE[39] = 11; assign amogusRLE[40] = 1; assign amogusRLE[41] = 1; assign amogusRLE[42] = 1; assign amogusRLE[43] = 1; assign amogusRLE[44] = 1; assign amogusRLE[45] = 3; assign amogusRLE[46] = 1; assign amogusRLE[47] = 1; assign amogusRLE[48] = 1; assign amogusRLE[49] = 1; assign amogusRLE[50] = 1; assign amogusRLE[51] = 1; assign amogusRLE[52] = 1; assign amogusRLE[53] = 1; assign amogusRLE[54] = 2; assign amogusRLE[55] = 1; assign amogusRLE[56] = 1; assign amogusRLE[57] = 1; assign amogusRLE[58] = 1; assign amogusRLE[59] = 1; assign amogusRLE[60] = 3; assign amogusRLE[61] = 9; assign amogusRLE[62] = 3; assign amogusRLE[63] = 1; assign amogusRLE[64] = 1; assign amogusRLE[65] = 3; assign amogusRLE[66] = 1; assign amogusRLE[67] = 1; assign amogusRLE[68] = 1; assign amogusRLE[69] = 1; assign amogusRLE[70] = 1; assign amogusRLE[71] = 1; assign amogusRLE[72] = 1; assign amogusRLE[73] = 2; assign amogusRLE[74] = 1; assign amogusRLE[75] = 1; assign amogusRLE[76] = 1; assign amogusRLE[77] = 1; assign amogusRLE[78] = 1; assign amogusRLE[79] = 3; assign amogusRLE[80] = 1; assign amogusRLE[81] = 9; assign amogusRLE[82] = 1; assign amogusRLE[83] = 1; assign amogusRLE[84] = 1; assign amogusRLE[85] = 1; assign amogusRLE[86] = 1; assign amogusRLE[87] = 3; assign amogusRLE[88] = 1; assign amogusRLE[89] = 2; assign amogusRLE[90] = 1; assign amogusRLE[91] = 3; assign amogusRLE[92] = 2; assign amogusRLE[93] = 2; assign amogusRLE[94] = 3; assign amogusRLE[95] = 1; assign amogusRLE[96] = 3; assign amogusRLE[97] = 91; assign amogusRLE[98] = 10; assign amogusRLE[99] = 24; assign amogusRLE[100] = 2; assign amogusRLE[101] = 7; assign amogusRLE[102] = 4; assign amogusRLE[103] = 21; assign amogusRLE[104] = 2; assign amogusRLE[105] = 11; assign amogusRLE[106] = 2; assign amogusRLE[107] = 20; assign amogusRLE[108] = 1; assign amogusRLE[109] = 13; assign amogusRLE[110] = 2; assign amogusRLE[111] = 18; assign amogusRLE[112] = 2; assign amogusRLE[113] = 14; assign amogusRLE[114] = 1; assign amogusRLE[115] = 18; assign amogusRLE[116] = 2; assign amogusRLE[117] = 2; assign amogusRLE[118] = 9; assign amogusRLE[119] = 3; assign amogusRLE[120] = 2; assign amogusRLE[121] = 17; assign amogusRLE[122] = 1; assign amogusRLE[123] = 2; assign amogusRLE[124] = 2; assign amogusRLE[125] = 7; assign amogusRLE[126] = 2; assign amogusRLE[127] = 3; assign amogusRLE[128] = 1; assign amogusRLE[129] = 16; assign amogusRLE[130] = 2; assign amogusRLE[131] = 2; assign amogusRLE[132] = 1; assign amogusRLE[133] = 9; assign amogusRLE[134] = 1; assign amogusRLE[135] = 3; assign amogusRLE[136] = 1; assign amogusRLE[137] = 16; assign amogusRLE[138] = 2; assign amogusRLE[139] = 2; assign amogusRLE[140] = 2; assign amogusRLE[141] = 7; assign amogusRLE[142] = 2; assign amogusRLE[143] = 3; assign amogusRLE[144] = 2; assign amogusRLE[145] = 15; assign amogusRLE[146] = 1; assign amogusRLE[147] = 4; assign amogusRLE[148] = 9; assign amogusRLE[149] = 5; assign amogusRLE[150] = 1; assign amogusRLE[151] = 14; assign amogusRLE[152] = 2; assign amogusRLE[153] = 6; assign amogusRLE[154] = 4; assign amogusRLE[155] = 8; assign amogusRLE[156] = 1; assign amogusRLE[157] = 14; assign amogusRLE[158] = 2; assign amogusRLE[159] = 18; assign amogusRLE[160] = 1; assign amogusRLE[161] = 14; assign amogusRLE[162] = 1; assign amogusRLE[163] = 19; assign amogusRLE[164] = 1; assign amogusRLE[165] = 14; assign amogusRLE[166] = 1; assign amogusRLE[167] = 19; assign amogusRLE[168] = 1; assign amogusRLE[169] = 14; assign amogusRLE[170] = 1; assign amogusRLE[171] = 19; assign amogusRLE[172] = 1; assign amogusRLE[173] = 14; assign amogusRLE[174] = 1; assign amogusRLE[175] = 19; assign amogusRLE[176] = 2; assign amogusRLE[177] = 12; assign amogusRLE[178] = 1; assign amogusRLE[179] = 20; assign amogusRLE[180] = 2; assign amogusRLE[181] = 12; assign amogusRLE[182] = 1; assign amogusRLE[183] = 21; assign amogusRLE[184] = 1; assign amogusRLE[185] = 12; assign amogusRLE[186] = 1; assign amogusRLE[187] = 21; assign amogusRLE[188] = 1; assign amogusRLE[189] = 12; assign amogusRLE[190] = 1; assign amogusRLE[191] = 21; assign amogusRLE[192] = 1; assign amogusRLE[193] = 12; assign amogusRLE[194] = 1; assign amogusRLE[195] = 21; assign amogusRLE[196] = 1; assign amogusRLE[197] = 11; assign amogusRLE[198] = 2; assign amogusRLE[199] = 21; assign amogusRLE[200] = 1; assign amogusRLE[201] = 11; assign amogusRLE[202] = 1; assign amogusRLE[203] = 22; assign amogusRLE[204] = 1; assign amogusRLE[205] = 11; assign amogusRLE[206] = 1; assign amogusRLE[207] = 22; assign amogusRLE[208] = 1; assign amogusRLE[209] = 11; assign amogusRLE[210] = 1; assign amogusRLE[211] = 5; assign amogusRLE[212] = 9; assign amogusRLE[213] = 8; assign amogusRLE[214] = 1; assign amogusRLE[215] = 11; assign amogusRLE[216] = 1; assign amogusRLE[217] = 4; assign amogusRLE[218] = 1; assign amogusRLE[219] = 8; assign amogusRLE[220] = 2; assign amogusRLE[221] = 7; assign amogusRLE[222] = 1; assign amogusRLE[223] = 10; assign amogusRLE[224] = 2; assign amogusRLE[225] = 4; assign amogusRLE[226] = 1; assign amogusRLE[227] = 9; assign amogusRLE[228] = 1; assign amogusRLE[229] = 7; assign amogusRLE[230] = 1; assign amogusRLE[231] = 10; assign amogusRLE[232] = 2; assign amogusRLE[233] = 4; assign amogusRLE[234] = 1; assign amogusRLE[235] = 9; assign amogusRLE[236] = 1; assign amogusRLE[237] = 7; assign amogusRLE[238] = 1; assign amogusRLE[239] = 5; assign amogusRLE[240] = 6; assign amogusRLE[241] = 6; assign amogusRLE[242] = 1; assign amogusRLE[243] = 8; assign amogusRLE[244] = 1; assign amogusRLE[245] = 7; assign amogusRLE[246] = 1; assign amogusRLE[247] = 4; assign amogusRLE[248] = 2; assign amogusRLE[249] = 4; assign amogusRLE[250] = 1; assign amogusRLE[251] = 6; assign amogusRLE[252] = 1; assign amogusRLE[253] = 8; assign amogusRLE[254] = 1; assign amogusRLE[255] = 7; assign amogusRLE[256] = 1; assign amogusRLE[257] = 4; assign amogusRLE[258] = 1; assign amogusRLE[259] = 12; assign amogusRLE[260] = 1; assign amogusRLE[261] = 7; assign amogusRLE[262] = 2; assign amogusRLE[263] = 7; assign amogusRLE[264] = 1; assign amogusRLE[265] = 4; assign amogusRLE[266] = 1; assign amogusRLE[267] = 11; assign amogusRLE[268] = 2; assign amogusRLE[269] = 4; assign amogusRLE[270] = 4; assign amogusRLE[271] = 8; assign amogusRLE[272] = 1; assign amogusRLE[273] = 5; assign amogusRLE[274] = 2; assign amogusRLE[275] = 7; assign amogusRLE[276] = 3; assign amogusRLE[277] = 4; assign amogusRLE[278] = 2; assign amogusRLE[279] = 11; assign amogusRLE[280] = 1; assign amogusRLE[281] = 6; assign amogusRLE[282] = 9; assign amogusRLE[283] = 5; assign amogusRLE[284] = 2; assign amogusRLE[285] = 12; assign amogusRLE[286] = 1; assign amogusRLE[287] = 20; assign amogusRLE[288] = 1; assign amogusRLE[289] = 12; assign amogusRLE[290] = 1; assign amogusRLE[291] = 21; assign amogusRLE[292] = 2; assign amogusRLE[293] = 9; assign amogusRLE[294] = 2; assign amogusRLE[295] = 24; assign amogusRLE[296] = 10; assign amogusRLE[297] = 28; assign amogusRLE[298] = 3; assign amogusRLE[299] = 44; assign amogusRLE[300] = 35;

  always @(posedge clk) begin
    if (reset) begin
      rle_segment_counter <= 0;
      rle_pixel_counter   <= 0;
      rle_pixel_state     <= start_pixel;

      line_pixel_counter  <= 0;
    end else begin
      rle_segment_counter <= next_rle_segment_counter;
      rle_pixel_counter <= next_rle_pixel_counter;
      rle_pixel_state <= next_rle_pixel_state;

      line_pixel_counter <= next_line_pixel_counter;
    end
  end

  always @(*) begin
    next_rle_segment_counter = rle_segment_counter;
    next_rle_pixel_counter = rle_pixel_counter;
    next_rle_pixel_state = rle_pixel_state;

    next_line_pixel_counter = line_pixel_counter;

    //default, if(img_sel == 0) begin
    current_rle_length     = logoRLE[rle_segment_counter];
    current_rle_n_segments = LEN_logoRLE;
    start_pixel = START_logoRLE;
    img_width = WIDTH_logoRLE;

    if(img_sel == 0) begin
      current_rle_length     = lambdaRLE[rle_segment_counter];
      current_rle_n_segments = LEN_lambdaRLE;
      start_pixel = START_lambdaRLE;
      img_width = WIDTH_lambdaRLE;
    end else if(img_sel == 2) begin
      current_rle_length     = intRLE[rle_segment_counter];
      current_rle_n_segments = LEN_intRLE;
      start_pixel = START_intRLE;
      img_width = WIDTH_intRLE;
    end
    /*
    else if(img_sel == 3) begin
      current_rle_length     = amogusRLE[rle_segment_counter];
      current_rle_n_segments = LEN_amogusRLE;
      start_pixel = START_amogusRLE;
      img_width = WIDTH_amogusRLE;
    end
    */
    
    
    h_sync = (line_pixel_counter == 0);
    v_sync = (rle_segment_counter == 0) && (rle_pixel_counter == 0);
    
    if(line_pixel_counter < img_width-1) begin
      next_line_pixel_counter = line_pixel_counter + 1;
    end else begin
      next_line_pixel_counter = 0;
    end
    
    if(rle_pixel_counter < current_rle_length-1) begin
      next_rle_pixel_counter = rle_pixel_counter + 1;
    end else begin
      next_rle_pixel_counter = 0;
      next_rle_pixel_state = !rle_pixel_state;

      if(rle_segment_counter < current_rle_n_segments-1) begin
        next_rle_segment_counter = rle_segment_counter + 1;
      end else begin
        next_rle_segment_counter = 0;
        next_rle_pixel_state = start_pixel;
        next_line_pixel_counter = 0;
      end
    end



    tx_out = enable_horizontal & ((line_pixel_counter == 0) | (line_pixel_counter == (img_width-1)));
    tx_out = tx_out | rle_pixel_state;
  end


endmodule