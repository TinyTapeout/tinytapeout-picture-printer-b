`timescale 1ns / 1ps
//`include "user_module_341542971476279892.v"

module user_module_341542971476279892_tb;



endmodule
